//Specification
package Spec;

parameter INST_LENGTH = 31;

typedef bit [INST_LENGTH:0] Instruction;

endpackage
