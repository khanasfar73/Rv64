//Specification
package Spec;

parameter INST_LENGTH = 63;

typedef bit [INST_LENGTH:0] Instruction;

endpackage
